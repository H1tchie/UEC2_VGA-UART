/**
 *  Copyright (C) 2023  AGH University of Science and Technology
 * MTM UEC2
 * Author: Piotr Kaczmarczyk
 *
 * Description:
 * Testbench for vga_timing module.
 */

`timescale 1 ns / 1 ps

module vga_timing_tb;

import vga_pkg::*;


/**
 *  Local parameters
 */

localparam CLK_PERIOD = 25;     // 40 MHz


/**
 * Local variables and signals
 */

logic clk;
logic rst;

wire [10:0] vcount, hcount;
wire        vsync,  hsync;
wire        vblnk,  hblnk;


/**
 * Clock generation
 */

initial begin
    clk = 1'b0;
    forever #(CLK_PERIOD/2) clk = ~clk;
end


/**
 * Reset generation
 */

initial begin
                       rst = 1'b0;
    #(1.25*CLK_PERIOD) rst = 1'b1;
                       rst = 1'b1;
    #(2.00*CLK_PERIOD) rst = 1'b0;
    zero();
end


/**
 * Dut placement
 */

vga_timing dut(
    .clk,
    .rst,
    .vcount,
    .vsync,
    .vblnk,
    .hcount,
    .hsync,
    .hblnk
);

/**
 * Tasks and functions
 */

 // Here you can declare tasks with immediate assertions (assert).
 
 task zero;
 
assert (hcount == 0 && vcount == 0)// $display ("We are at the top left corner of screen");
     else $error("reset nie dziala");
 

endtask
/**
 */

// Here you can declare concurrent assertions (assert property).

 // UWAGA 2 PIERWSZE ERRORY Z KAZDEJ ASSERCJI WYNIKAJA Z STANU NIEUSTALONEGO NA POCZATKU SYMULACJI
// NIEBRAC ICH POD UWAGE PRZY DEBUGOWANIU
 assert property (@(posedge clk)hcount<=HOR_MAX || hcount === 'x )// $display ("hcoount jest w zakresie");
    else $error("hcount poza zakresem");
assert property (@(posedge clk)vcount<=VER_MAX ||vcount === 'x)// $display ("vcount jest w zakresie");
    else $error("vcount poza zakresem");
assert property (@(posedge clk)((vcount > VER_SYNCH_START-1) && (vcount < VER_SYNCH_STOP) & vsync == 1) || vcount === 'x|| ((vcount <= VER_SYNCH_START-1) || (vcount >= VER_SYNCH_STOP) & vsync == 0) )
    else $error("synchronizacja wertykalna nie dziala");
assert property (@(posedge clk)((hcount > HOR_SYNCH_START-1) && (hcount < HOR_SYNCH_STOP) & hsync == 1) || hcount === 'x|| ((hcount <= HOR_SYNCH_START-1) || (hcount >= HOR_SYNCH_STOP) & hsync == 0) )
    else $error("synchronizacja horyzontalna nie dziala");
assert property (@(posedge clk)(vcount>= VER_BLANK_START && vblnk == 1)|| vcount === 'x||(vcount<VER_BLANK_START && vblnk == 0))
    else $error("blanking wertykalny nie dziala");
assert property (@(posedge clk)(hcount>= HOR_BLANK_START && hblnk == 1)||hcount === 'x||(hcount<HOR_BLANK_START && hblnk == 0))
    else $error("blanking horyzontalny nie dziala");


/**
 * Main test
 */

initial begin
    @(posedge rst);
    @(negedge rst);

    wait (vsync == 1'b0);
    @(negedge vsync)
    @(negedge vsync)

    $finish;
end

endmodule
